// Automatisch generierte Defines aus .config Datei
// NICHT MANUELL BEARBEITEN!
// Generiert am: 2025-09-24 14:31:06

`define FILTER_SIZE 3
`define DATA_WIDTH 8
`define IMAGE_CHANNELS 1
`define IMAGE_PATCH_SIZE 3

// Parameter als SystemVerilog Parameter
parameter int FILTER_SIZE = `FILTER_SIZE;
parameter int DATA_WIDTH = `DATA_WIDTH;
parameter int IMAGE_CHANNELS = `IMAGE_CHANNELS;
parameter int IMAGE_PATCH_SIZE = `IMAGE_PATCH_SIZE;
